LIBRARY IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;
entity InstrMem32bit is
	port (
	        address  : in STD_LOGIC_VECTOR (31 downto 0);
		      Instr    : out STD_LOGIC_VECTOR (31 downto 0)
		    );
end InstrMem32bit;

architecture Behavioral of InstrMem32bit is
	Type rom_type is ARRAY (0 to 255) of STD_LOGIC_VECTOR(31 downto 0);
	Signal Rom : rom_type := (	X"2000000F",X"20210002",X"20420001",X"20630001",X"20c60000",X"20c60000",X"aca20000",X"aca30001",X"20210001",X"20420001",X"20630002",X"20c60000",X"20210001",X"aca20000",X"aca30001",X"20c60000",X"20210001",X"20420003",X"20630005",X"20c60000",X"20210001",X"aca20000",X"aca30001",X"20c60000",X"20210001",X"20420008",X"2063000d",X"20c60000",X"20210001",X"aca20000",X"aca30001"
	,X"20c60000",X"20210001",X"20420015",X"20630022",X"20c60000",X"20210001",X"aca20000",X"aca30001",X"20c60000",X"20210001",X"20420037",X"20630059",X"20c60000",X"20210001",X"aca20000",X"aca30001"
	,X"20c60000",X"20210001",X"20420090",X"206300e9",X"20c60000",X"20210001",X"aca20000",X"aca30001",X"20c60000",X"20210001",X"20420179",X"20630000",X"20c60000",X"20210000",X"aca20000",X"aca30001",X"00000000",X"00000000",
											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"	);											
	begin
		Instr <= Rom ( to_integer(unsigned(address)));
end Behavioral;